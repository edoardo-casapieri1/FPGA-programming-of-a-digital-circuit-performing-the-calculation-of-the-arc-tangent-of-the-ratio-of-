library IEEE; 
use IEEE.std_logic_1164.all;

entity Cordic_tb is
end entity Cordic_tb;

architecture test of Cordic_tb is

constant T_CLK: time := 12 ns;
constant N_tb : integer := 12;

signal clk_tb : std_logic := '0';
signal end_sim : std_logic := '0';

signal ready_tb : std_logic := '0';  
						      
signal ingr_x_tb : std_logic_vector (11 downto 0) := "000000000010"; -- Inserire qui il valore del denominatore
signal ingr_y_tb : std_logic_vector (11 downto 0) := "111111111110"; -- Inserire qui il valore del numeratore       
signal ris_tb : std_logic_vector(N_tb-1 downto 0);
          
component Cordic is
generic ( N : positive := 12);
   port( 
         cordic_den     :  in std_logic_VECTOR (11 downto 0);
         cordic_num     :  in std_logic_VECTOR (11 downto 0);
         cordic_ris       :  out std_logic_VECTOR (11 downto 0);
         cordic_clock          :  in  std_logic;
         cordic_ready       :  in  std_logic
    );
end component Cordic;

begin

    clk_tb <= not(clk_tb) or end_sim after T_CLK/2;
    ready_tb <= '1' after T_CLK, '0' after 3*T_CLK;
    end_sim <= '1' after 100*T_CLK;

    dut: CORDIC
    generic map (N => N_tb)
    port map(
                cordic_den => ingr_x_tb,
                cordic_num => ingr_y_tb,
                cordic_ris => ris_tb,
                cordic_clock => clk_tb,
                cordic_ready => ready_tb
    );
    
end architecture test;